-- ***** BEGIN LICENSE BLOCK *****
-- 
-- $Id: Divider.vhd,v 1.2 2006-10-05 16:17:11 petebleackley Exp $ $Name: not supported by cvs2svn $
-- *
-- * Version: MPL 1.1/GPL 2.0/LGPL 2.1
-- *
-- * The contents of this file are subject to the Mozilla Public License
-- * Version 1.1 (the "License"); you may not use this file except in compliance
-- * with the License. You may obtain a copy of the License at
-- * http://www.mozilla.org/MPL/
-- *
-- * Software distributed under the License is distributed on an "AS IS" basis,
-- * WITHOUT WARRANTY OF ANY KIND, either express or implied. See the License for
-- * the specific language governing rights and limitations under the License.
-- *
-- * The Original Code is BBC Research and Development code.
-- *
-- * The Initial Developer of the Original Code is the British Broadcasting
-- * Corporation.
-- * Portions created by the Initial Developer are Copyright (C) 2004.
-- * All Rights Reserved.
-- *
-- * Contributor(s): Peter Bleackley (Original author)
-- *
-- * Alternatively, the contents of this file may be used under the terms of
-- * the GNU General Public License Version 2 (the "GPL"), or the GNU Lesser
-- * Public License Version 2.1 (the "LGPL"), in which case the provisions of
-- * the GPL or the LGPL are applicable instead of those above. If you wish to
-- * allow use of your version of this file only under the terms of the either
-- * the GPL or LGPL and not to allow others to use your version of this file
-- * under the MPL, indicate your decision by deleting the provisions above
-- * and replace them with the notice and other provisions required by the GPL
-- * or LGPL. If you do not delete the provisions above, a recipient may use
-- * your version of this file under the terms of any one of the MPL, the GPL
-- * or the LGPL.
-- * ***** END LICENSE BLOCK ***** */

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

--  Uncomment the following lines to use the declarations that are
--  provided for instantiating Xilinx primitive components.
--library UNISIM;
--use UNISIM.VComponents.all;

entity Divider is
    Port ( NUMERATOR : in std_logic_vector(7 downto 0);
           DENOMINATOR : in std_logic_vector(7 downto 0);
			  RESET : in std_logic;
           CLOCK : in std_logic;
           QUOTIENT : out std_logic_vector(7 downto 0));
end Divider;

architecture RTL of Divider is
	signal NUMERATOR2 : std_logic_vector(7 downto 0);
	signal DENOMINATOR2 : std_logic_vector(7 downto 0);
	signal RECIPROCAL : std_logic_vector(15 downto 0);
	signal PRODUCT : std_logic_vector(23 downto 0);
	signal INDEX : std_logic_vector (7 downto 0);
	type ROM is array (253 downto 0) of std_logic_vector(15 downto 0);
	constant LUT : ROM :=  ( "0000000100000001",
"0000000100000010",
"0000000100000011",
"0000000100000100",
"0000000100000101",
"0000000100000110",
"0000000100000111",
"0000000100001000",
"0000000100001001",
"0000000100001010",
"0000000100001011",
"0000000100001101",
"0000000100001110",
"0000000100001111",
"0000000100010000",
"0000000100010001",
"0000000100010010",
"0000000100010011",
"0000000100010101",
"0000000100010110",
"0000000100010111",
"0000000100011000",
"0000000100011001",
"0000000100011010",
"0000000100011100",
"0000000100011101",
"0000000100011110",
"0000000100011111",
"0000000100100001",
"0000000100100010",
"0000000100100011",
"0000000100100101",
"0000000100100110",
"0000000100100111",
"0000000100101001",
"0000000100101010",
"0000000100101011",
"0000000100101101",
"0000000100101110",
"0000000100101111",
"0000000100110001",
"0000000100110010",
"0000000100110100",
"0000000100110101",
"0000000100110111",
"0000000100111000",
"0000000100111010",
"0000000100111011",
"0000000100111101",
"0000000100111110",
"0000000101000000",
"0000000101000001",
"0000000101000011",
"0000000101000100",
"0000000101000110",
"0000000101001000",
"0000000101001001",
"0000000101001011",
"0000000101001101",
"0000000101001110",
"0000000101010000",
"0000000101010010",
"0000000101010100",
"0000000101010101",
"0000000101010111",
"0000000101011001",
"0000000101011011",
"0000000101011101",
"0000000101011110",
"0000000101100000",
"0000000101100010",
"0000000101100100",
"0000000101100110",
"0000000101101000",
"0000000101101010",
"0000000101101100",
"0000000101101110",
"0000000101110000",
"0000000101110010",
"0000000101110100",
"0000000101110110",
"0000000101111001",
"0000000101111011",
"0000000101111101",
"0000000101111111",
"0000000110000010",
"0000000110000100",
"0000000110000110",
"0000000110001000",
"0000000110001011",
"0000000110001101",
"0000000110010000",
"0000000110010010",
"0000000110010101",
"0000000110010111",
"0000000110011010",
"0000000110011100",
"0000000110011111",
"0000000110100001",
"0000000110100100",
"0000000110100111",
"0000000110101010",
"0000000110101100",
"0000000110101111",
"0000000110110010",
"0000000110110101",
"0000000110111000",
"0000000110111011",
"0000000110111110",
"0000000111000001",
"0000000111000100",
"0000000111000111",
"0000000111001010",
"0000000111001110",
"0000000111010001",
"0000000111010100",
"0000000111010111",
"0000000111011011",
"0000000111011110",
"0000000111100010",
"0000000111100101",
"0000000111101001",
"0000000111101101",
"0000000111110000",
"0000000111110100",
"0000000111111000",
"0000000111111100",
"0000001000000000",
"0000001000000100",
"0000001000001000",
"0000001000001100",
"0000001000010001",
"0000001000010101",
"0000001000011001",
"0000001000011110",
"0000001000100010",
"0000001000100111",
"0000001000101011",
"0000001000110000",
"0000001000110101",
"0000001000111010",
"0000001000111111",
"0000001001000100",
"0000001001001001",
"0000001001001110",
"0000001001010100",
"0000001001011001",
"0000001001011111",
"0000001001100100",
"0000001001101010",
"0000001001110000",
"0000001001110110",
"0000001001111100",
"0000001010000011",
"0000001010001001",
"0000001010001111",
"0000001010010110",
"0000001010011101",
"0000001010100100",
"0000001010101011",
"0000001010110010",
"0000001010111001",
"0000001011000001",
"0000001011001000",
"0000001011010000",
"0000001011011000",
"0000001011100000",
"0000001011101001",
"0000001011110001",
"0000001011111010",
"0000001100000011",
"0000001100001100",
"0000001100010110",
"0000001100011111",
"0000001100101001",
"0000001100110011",
"0000001100111110",
"0000001101001000",
"0000001101010011",
"0000001101011110",
"0000001101101010",
"0000001101110110",
"0000001110000010",
"0000001110001110",
"0000001110011011",
"0000001110101000",
"0000001110110110",
"0000001111000100",
"0000001111010010",
"0000001111100001",
"0000001111110000",
"0000010000000000",
"0000010000010000",
"0000010000100001",
"0000010000110010",
"0000010001000100",
"0000010001010111",
"0000010001101010",
"0000010001111110",
"0000010010010010",
"0000010010101000",
"0000010010111110",
"0000010011010101",
"0000010011101100",
"0000010100000101",
"0000010100011111",
"0000010100111001",
"0000010101010101",
"0000010101110010",
"0000010110010001",
"0000010110110000",
"0000010111010001",
"0000010111110100",
"0000011000011000",
"0000011000111110",
"0000011001100110",
"0000011010010000",
"0000011010111101",
"0000011011101011",
"0000011100011100",
"0000011101010000",
"0000011110001000",
"0000011111000010",
"0000100000000000",
"0000100001000010",
"0000100010001001",
"0000100011010100",
"0000100100100101",
"0000100101111011",
"0000100111011001",
"0000101000111101",
"0000101010101011",
"0000101100100001",
"0000101110100011",
"0000110000110001",
"0000110011001101",
"0000110101111001",
"0000111000111001",
"0000111100001111",
"0001000000000000",
"0001000100010001",
"0001001001001001",
"0001001110110001",
"0001010101010101",
"0001011101000110",
"0001100110011010",
"0001110001110010",
"0010000000000000",
"0010010010010010",
"0010101010101011",
"0011001100110011",
"0100000000000000",
"0101010101010101",
"1000000000000000");
begin

INIT : process(DENOMINATOR,RESET)
begin
	if RESET = '1' then
		DENOMINATOR2 <= "00000010";
	else
		DENOMINATOR2 <= DENOMINATOR;
	end if;
end process INIT;

SETNUMERATOR : process (CLOCK)
begin
	if CLOCK'event and CLOCK = '1' then
		if RESET = '1' then
			NUMERATOR2 <= "00000001";
		else
			NUMERATOR2 <= NUMERATOR;
		end if;
	end if;
end process SETNUMERATOR;
			

INDEX <= DENOMINATOR2 - "00000010";

LOOKUP: process(CLOCK)
begin
	if CLOCK'event and CLOCK = '1' then
		 RECIPROCAL <= LUT(conv_integer(INDEX));
	end if;
end process LOOKUP;

DIVIDE: process(CLOCK)
begin
	if CLOCK'event and CLOCK='1' then
		PRODUCT<=NUMERATOR2*RECIPROCAL;
	end if;
end process DIVIDE;


QUOTIENT <=	 PRODUCT(15 downto 8);


end RTL;
