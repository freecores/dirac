-- ***** BEGIN LICENSE BLOCK *****
-- 
-- 
--  Version: MPL 1.1/GPL 2.0/LGPL 2.1
-- 
--  The contents of this file are subject to the Mozilla Public License
--  Version 1.1 (the "License"); you may not use this file except in compliance
--  with the License. You may obtain a copy of the License at
--  http://www.mozilla.org/MPL/
-- 
--  Software distributed under the License is distributed on an "AS IS" basis,
--  WITHOUT WARRANTY OF ANY KIND, either express or implied. See the License for
--  the specific language governing rights and limitations under the License.
-- 
--  The Original Code is BBC Research and Development code.
-- 
--  The Initial Developer of the Original Code is the British Broadcasting
--  Corporation.
--  Portions created by the Initial Developer are Copyright (C) 2006.
--  All Rights Reserved.
-- 
--  Contributor(s): Peter Bleackley (Original author)
-- 
--  Alternatively, the contents of this file may be used under the terms of
--  the GNU General Public License Version 2 (the "GPL"), or the GNU Lesser
--  Public License Version 2.1 (the "LGPL"), in which case the provisions of
--  the GPL or the LGPL are applicable instead of those above. If you wish to
--  allow use of your version of this file only under the terms of the either
--  the GPL or LGPL and not to allow others to use your version of this file
--  under the MPL, indicate your decision by deleting the provisions above
--  and replace them with the notice and other provisions required by the GPL
--  or LGPL. If you do not delete the provisions above, a recipient may use
--  your version of this file under the terms of any one of the MPL, the GPL
--  or the LGPL.
-- * ***** END LICENSE BLOCK ***** */

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

--  Uncomment the following lines to use the declarations that are
--  provided for instantiating Xilinx primitive components.
--library UNISIM;
--use UNISIM.VComponents.all;

entity Divider is
    Port ( NUMERATOR : in std_logic_vector(9 downto 0);
           DENOMINATOR : in std_logic_vector(9 downto 0);
			  RESET : in std_logic;
           CLOCK : in std_logic;
           QUOTIENT : out std_logic_vector(9 downto 0));
end Divider;

architecture RTL of Divider is
	signal NUMERATOR2 : std_logic_vector(9 downto 0);
	signal DENOMINATOR2 : std_logic_vector( 9 downto 0);
	signal RECIPROCAL : std_logic_vector(31 downto 0);
	signal PRODUCT1 : std_logic_vector(25 downto 0);
	signal PRODUCT2 : std_logic_vector(25 downto 0);
	signal TOTAL : std_logic_vector(41 downto 0);
	signal INDEX : std_logic_vector (9 downto 0);
	type ROM is array (1021 downto 0) of std_logic_vector(31 downto 0);
	constant LUT : ROM :=  ("00000000010000000001000000000100",
"00000000010000000010000000010000",
"00000000010000000011000000100100",
"00000000010000000100000001000000",
"00000000010000000101000001100100",
"00000000010000000110000010010000",
"00000000010000000111000011000101",
"00000000010000001000000100000010",
"00000000010000001001000101000110",
"00000000010000001010000110010011",
"00000000010000001011000111101001",
"00000000010000001100001001000110",
"00000000010000001101001010101100",
"00000000010000001110001100011010",
"00000000010000001111001110010001",
"00000000010000010000010000010000",
"00000000010000010001010010010111",
"00000000010000010010010100100111",
"00000000010000010011010110111111",
"00000000010000010100011001011111",
"00000000010000010101011100001000",
"00000000010000010110011110111010",
"00000000010000010111100001110100",
"00000000010000011000100100110111",
"00000000010000011001101000000010",
"00000000010000011010101011010110",
"00000000010000011011101110110010",
"00000000010000011100110010011000",
"00000000010000011101110110000110",
"00000000010000011110111001111100",
"00000000010000011111111101111100",
"00000000010000100001000010000100",
"00000000010000100010000110010101",
"00000000010000100011001010101110",
"00000000010000100100001111010001",
"00000000010000100101010011111100",
"00000000010000100110011000110001",
"00000000010000100111011101101110",
"00000000010000101000100010110100",
"00000000010000101001101000000100",
"00000000010000101010101101011100",
"00000000010000101011110010111101",
"00000000010000101100111000101000",
"00000000010000101101111110011011",
"00000000010000101111000100011000",
"00000000010000110000001010011110",
"00000000010000110001010000101101",
"00000000010000110010010111000101",
"00000000010000110011011101100110",
"00000000010000110100100100010001",
"00000000010000110101101011000101",
"00000000010000110110110010000010",
"00000000010000110111111001001001",
"00000000010000111001000000011001",
"00000000010000111010000111110010",
"00000000010000111011001111010101",
"00000000010000111100010111000010",
"00000000010000111101011110110111",
"00000000010000111110100110110111",
"00000000010000111111101111000000",
"00000000010001000000110111010010",
"00000000010001000001111111101110",
"00000000010001000011001000010100",
"00000000010001000100010001000100",
"00000000010001000101011001111101",
"00000000010001000110100011000000",
"00000000010001000111101100001101",
"00000000010001001000110101100011",
"00000000010001001001111111000011",
"00000000010001001011001000101110",
"00000000010001001100010010100010",
"00000000010001001101011100100000",
"00000000010001001110100110101000",
"00000000010001001111110000111010",
"00000000010001010000111011010110",
"00000000010001010010000101111100",
"00000000010001010011010000101100",
"00000000010001010100011011100110",
"00000000010001010101100110101010",
"00000000010001010110110001111001",
"00000000010001010111111101010010",
"00000000010001011001001000110101",
"00000000010001011010010100100010",
"00000000010001011011100000011010",
"00000000010001011100101100011100",
"00000000010001011101111000101000",
"00000000010001011111000100111111",
"00000000010001100000010001100000",
"00000000010001100001011110001011",
"00000000010001100010101011000010",
"00000000010001100011111000000010",
"00000000010001100101000101001110",
"00000000010001100110010010100011",
"00000000010001100111100000000100",
"00000000010001101000101101101111",
"00000000010001101001111011100101",
"00000000010001101011001001100110",
"00000000010001101100010111110001",
"00000000010001101101100110000111",
"00000000010001101110110100101001",
"00000000010001110000000011010101",
"00000000010001110001010010001011",
"00000000010001110010100001001101",
"00000000010001110011110000011010",
"00000000010001110100111111110010",
"00000000010001110110001111010101",
"00000000010001110111011111000011",
"00000000010001111000101110111100",
"00000000010001111001111111000001",
"00000000010001111011001111010000",
"00000000010001111100011111101011",
"00000000010001111101110000010001",
"00000000010001111111000001000011",
"00000000010010000000010010000000",
"00000000010010000001100011001000",
"00000000010010000010110100011100",
"00000000010010000100000101111011",
"00000000010010000101010111100110",
"00000000010010000110101001011100",
"00000000010010000111111011011110",
"00000000010010001001001101101011",
"00000000010010001010100000000100",
"00000000010010001011110010101001",
"00000000010010001101000101011001",
"00000000010010001110011000010110",
"00000000010010001111101011011110",
"00000000010010010000111110110010",
"00000000010010010010010010010010",
"00000000010010010011100101111110",
"00000000010010010100111001110101",
"00000000010010010110001101111001",
"00000000010010010111100010001001",
"00000000010010011000110110100101",
"00000000010010011010001011001101",
"00000000010010011011100000000010",
"00000000010010011100110101000010",
"00000000010010011110001010001111",
"00000000010010011111011111101000",
"00000000010010100000110101001110",
"00000000010010100010001011000000",
"00000000010010100011100000111110",
"00000000010010100100110111001001",
"00000000010010100110001101100000",
"00000000010010100111100100000100",
"00000000010010101000111010110101",
"00000000010010101010010001110010",
"00000000010010101011101000111100",
"00000000010010101101000000010010",
"00000000010010101110010111110110",
"00000000010010101111101111100110",
"00000000010010110001000111100011",
"00000000010010110010011111101101",
"00000000010010110011111000000100",
"00000000010010110101010000101000",
"00000000010010110110101001011000",
"00000000010010111000000010010111",
"00000000010010111001011011100010",
"00000000010010111010110100111010",
"00000000010010111100001110100000",
"00000000010010111101101000010010",
"00000000010010111111000010010011",
"00000000010011000000011100100000",
"00000000010011000001110110111011",
"00000000010011000011010001100100",
"00000000010011000100101100011001",
"00000000010011000110000111011101",
"00000000010011000111100010101110",
"00000000010011001000111110001101",
"00000000010011001010011001111001",
"00000000010011001011110101110011",
"00000000010011001101010001111011",
"00000000010011001110101110010001",
"00000000010011010000001010110101",
"00000000010011010001100111100110",
"00000000010011010011000100100110",
"00000000010011010100100001110011",
"00000000010011010101111111001111",
"00000000010011010111011100111001",
"00000000010011011000111010110001",
"00000000010011011010011000110111",
"00000000010011011011110111001100",
"00000000010011011101010101101111",
"00000000010011011110110100100000",
"00000000010011100000010011100000",
"00000000010011100001110010101110",
"00000000010011100011010010001011",
"00000000010011100100110001110110",
"00000000010011100110010001110000",
"00000000010011100111110001111001",
"00000000010011101001010010010000",
"00000000010011101010110010110111",
"00000000010011101100010011101100",
"00000000010011101101110100110000",
"00000000010011101111010110000011",
"00000000010011110000110111100101",
"00000000010011110010011001010110",
"00000000010011110011111011010110",
"00000000010011110101011101100110",
"00000000010011110111000000000100",
"00000000010011111000100010110010",
"00000000010011111010000101110000",
"00000000010011111011101000111101",
"00000000010011111101001100011001",
"00000000010011111110110000000100",
"00000000010100000000010100000000",
"00000000010100000001111000001011",
"00000000010100000011011100100101",
"00000000010100000101000001010000",
"00000000010100000110100110001010",
"00000000010100001000001011010100",
"00000000010100001001110000101110",
"00000000010100001011010110011000",
"00000000010100001100111100010010",
"00000000010100001110100010011100",
"00000000010100010000001000110111",
"00000000010100010001101111100001",
"00000000010100010011010110011100",
"00000000010100010100111101100111",
"00000000010100010110100101000011",
"00000000010100011000001100101111",
"00000000010100011001110100101011",
"00000000010100011011011100111000",
"00000000010100011101000101010110",
"00000000010100011110101110000101",
"00000000010100100000010111000100",
"00000000010100100010000000010100",
"00000000010100100011101001110101",
"00000000010100100101010011100111",
"00000000010100100110111101101010",
"00000000010100101000100111111110",
"00000000010100101010010010100011",
"00000000010100101011111101011010",
"00000000010100101101101000100010",
"00000000010100101111010011111011",
"00000000010100110000111111100110",
"00000000010100110010101011100010",
"00000000010100110100010111101111",
"00000000010100110110000100001110",
"00000000010100110111110000111111",
"00000000010100111001011110000010",
"00000000010100111011001011010111",
"00000000010100111100111000111101",
"00000000010100111110100110110101",
"00000000010101000000010101000000",
"00000000010101000010000011011100",
"00000000010101000011110010001011",
"00000000010101000101100001001100",
"00000000010101000111010000011111",
"00000000010101001001000000000101",
"00000000010101001010101111111101",
"00000000010101001100100000000111",
"00000000010101001110010000100101",
"00000000010101010000000001010101",
"00000000010101010001110010010111",
"00000000010101010011100011101101",
"00000000010101010101010101010101",
"00000000010101010111000111010000",
"00000000010101011000111001011110",
"00000000010101011010101100000000",
"00000000010101011100011110110100",
"00000000010101011110010001111100",
"00000000010101100000000101011000",
"00000000010101100001111001000110",
"00000000010101100011101101001000",
"00000000010101100101100001011110",
"00000000010101100111010110000111",
"00000000010101101001001011000100",
"00000000010101101011000000010101",
"00000000010101101100110101111010",
"00000000010101101110101011110011",
"00000000010101110000100001111111",
"00000000010101110010011000100000",
"00000000010101110100001111010101",
"00000000010101110110000110011111",
"00000000010101110111111101111100",
"00000000010101111001110101101110",
"00000000010101111011101101110101",
"00000000010101111101100110010000",
"00000000010101111111011111000000",
"00000000010110000001011000000101",
"00000000010110000011010001011111",
"00000000010110000101001011001101",
"00000000010110000111000101010001",
"00000000010110001000111111101001",
"00000000010110001010111010010111",
"00000000010110001100110101011010",
"00000000010110001110110000110011",
"00000000010110010000101100100001",
"00000000010110010010101000100100",
"00000000010110010100100100111110",
"00000000010110010110100001101100",
"00000000010110011000011110110001",
"00000000010110011010011100001100",
"00000000010110011100011001111100",
"00000000010110011110011000000011",
"00000000010110100000010110100000",
"00000000010110100010010101010011",
"00000000010110100100010100011100",
"00000000010110100110010011111100",
"00000000010110101000010011110011",
"00000000010110101010010100000000",
"00000000010110101100010100100100",
"00000000010110101110010101011110",
"00000000010110110000010110110000",
"00000000010110110010011000011000",
"00000000010110110100011010011000",
"00000000010110110110011100101111",
"00000000010110111000011111011101",
"00000000010110111010100010100011",
"00000000010110111100100110000000",
"00000000010110111110101001110101",
"00000000010111000000101110000001",
"00000000010111000010110010100101",
"00000000010111000100110111100001",
"00000000010111000110111100110101",
"00000000010111001001000010100001",
"00000000010111001011001000100110",
"00000000010111001101001111000011",
"00000000010111001111010101111000",
"00000000010111010001011101000101",
"00000000010111010011100100101100",
"00000000010111010101101100101011",
"00000000010111010111110101000010",
"00000000010111011001111101110011",
"00000000010111011100000110111101",
"00000000010111011110010000100000",
"00000000010111100000011010011100",
"00000000010111100010100100110010",
"00000000010111100100101111100001",
"00000000010111100110111010101001",
"00000000010111101001000110001100",
"00000000010111101011010010001000",
"00000000010111101101011110011110",
"00000000010111101111101011001110",
"00000000010111110001111000011000",
"00000000010111110100000101111101",
"00000000010111110110010011111011",
"00000000010111111000100010010101",
"00000000010111111010110001001001",
"00000000010111111101000000010111",
"00000000010111111111010000000001",
"00000000011000000001100000000110",
"00000000011000000011110000100101",
"00000000011000000110000001100000",
"00000000011000001000010010110110",
"00000000011000001010100100101000",
"00000000011000001100110110110101",
"00000000011000001111001001011101",
"00000000011000010001011100100010",
"00000000011000010011110000000011",
"00000000011000010110000011111111",
"00000000011000011000011000011000",
"00000000011000011010101101001101",
"00000000011000011101000010011110",
"00000000011000011111011000001101",
"00000000011000100001101110010111",
"00000000011000100100000100111111",
"00000000011000100110011100000011",
"00000000011000101000110011100101",
"00000000011000101011001011100100",
"00000000011000101101100100000000",
"00000000011000101111111100111010",
"00000000011000110010010110010001",
"00000000011000110100110000000110",
"00000000011000110111001010011001",
"00000000011000111001100101001001",
"00000000011000111100000000011000",
"00000000011000111110011100000110",
"00000000011001000000111000010001",
"00000000011001000011010100111100",
"00000000011001000101110010000101",
"00000000011001001000001111101101",
"00000000011001001010101101110100",
"00000000011001001101001100011001",
"00000000011001001111101011011111",
"00000000011001010010001011000011",
"00000000011001010100101011001000",
"00000000011001010111001011101100",
"00000000011001011001101100110000",
"00000000011001011100001110010011",
"00000000011001011110110000010111",
"00000000011001100001010010111100",
"00000000011001100011110110000000",
"00000000011001100110011001100110",
"00000000011001101000111101101100",
"00000000011001101011100010010011",
"00000000011001101110000111011011",
"00000000011001110000101101000101",
"00000000011001110011010011010000",
"00000000011001110101111001111100",
"00000000011001111000100001001010",
"00000000011001111011001000111010",
"00000000011001111101110001001100",
"00000000011010000000011010000000",
"00000000011010000011000011010110",
"00000000011010000101101101001111",
"00000000011010001000010111101011",
"00000000011010001011000010101010",
"00000000011010001101101110001011",
"00000000011010010000011010010000",
"00000000011010010011000110111000",
"00000000011010010101110100000100",
"00000000011010011000100001110011",
"00000000011010011011010000000110",
"00000000011010011101111110111101",
"00000000011010100000101110011001",
"00000000011010100011011110011001",
"00000000011010100110001110111101",
"00000000011010101001000000000110",
"00000000011010101011110001110100",
"00000000011010101110100100000111",
"00000000011010110001010111000000",
"00000000011010110100001010011110",
"00000000011010110110111110100001",
"00000000011010111001110011001011",
"00000000011010111100101000011010",
"00000000011010111111011110010000",
"00000000011011000010010100101100",
"00000000011011000101001011101111",
"00000000011011001000000011011001",
"00000000011011001010111011101001",
"00000000011011001101110100100001",
"00000000011011010000101110000000",
"00000000011011010011101000000110",
"00000000011011010110100010110101",
"00000000011011011001011110001011",
"00000000011011011100011010001010",
"00000000011011011111010110110000",
"00000000011011100010010100000000",
"00000000011011100101010001111000",
"00000000011011101000010000011001",
"00000000011011101011001111100100",
"00000000011011101110001111011000",
"00000000011011110001001111110101",
"00000000011011110100010000111100",
"00000000011011110111010010101110",
"00000000011011111010010101001001",
"00000000011011111101011000001111",
"00000000011100000000011100000000",
"00000000011100000011100000011100",
"00000000011100000110100101100010",
"00000000011100001001101011010100",
"00000000011100001100110001110010",
"00000000011100001111111000111100",
"00000000011100010011000000110001",
"00000000011100010110001001010011",
"00000000011100011001010010100001",
"00000000011100011100011100011100",
"00000000011100011111100111000100",
"00000000011100100010110010011001",
"00000000011100100101111110011011",
"00000000011100101001001011001100",
"00000000011100101100011000101010",
"00000000011100101111100110110110",
"00000000011100110010110101110000",
"00000000011100110110000101011010",
"00000000011100111001010101110010",
"00000000011100111100100110111001",
"00000000011100111111111000110000",
"00000000011101000011001011010110",
"00000000011101000110011110101100",
"00000000011101001001110010110010",
"00000000011101001101000111101001",
"00000000011101010000011101010000",
"00000000011101010011110011101000",
"00000000011101010111001010110010",
"00000000011101011010100010101100",
"00000000011101011101111011011001",
"00000000011101100001010100110111",
"00000000011101100100101111001000",
"00000000011101101000001010001011",
"00000000011101101011100110000001",
"00000000011101101111000010101010",
"00000000011101110010100000000111",
"00000000011101110101111110010111",
"00000000011101111001011101011011",
"00000000011101111100111101010011",
"00000000011110000000011110000000",
"00000000011110000011111111100001",
"00000000011110000111100001111000",
"00000000011110001011000101000100",
"00000000011110001110101001000101",
"00000000011110010010001101111101",
"00000000011110010101110011101011",
"00000000011110011001011010001111",
"00000000011110011101000001101010",
"00000000011110100000101001111100",
"00000000011110100100010011000110",
"00000000011110100111111101001000",
"00000000011110101011101000000001",
"00000000011110101111010011110011",
"00000000011110110011000000011110",
"00000000011110110110101110000010",
"00000000011110111010011100011111",
"00000000011110111110001011110110",
"00000000011111000001111100000111",
"00000000011111000101101101010011",
"00000000011111001001011111011001",
"00000000011111001101010010011010",
"00000000011111010001000110010110",
"00000000011111010100111011001110",
"00000000011111011000110001000010",
"00000000011111011100100111110011",
"00000000011111100000011111100000",
"00000000011111100100011000001010",
"00000000011111101000010001110010",
"00000000011111101100001100011000",
"00000000011111110000000111111100",
"00000000011111110100000100011110",
"00000000011111111000000001111111",
"00000000011111111100000000011111",
"00000000100000000000000000000000",
"00000000100000000100000000100000",
"00000000100000001000000010000000",
"00000000100000001100000100100001",
"00000000100000010000001000000100",
"00000000100000010100001100100111",
"00000000100000011000010010001101",
"00000000100000011100011000110101",
"00000000100000100000100000100000",
"00000000100000100100101001001110",
"00000000100000101000110010111111",
"00000000100000101100111101110101",
"00000000100000110001001001101110",
"00000000100000110101010110101100",
"00000000100000111001100100110000",
"00000000100000111101110011111001",
"00000000100001000010000100001000",
"00000000100001000110010101011101",
"00000000100001001010100111111001",
"00000000100001001110111011011101",
"00000000100001010011010000001000",
"00000000100001010111100101111011",
"00000000100001011011111100110111",
"00000000100001100000010100111100",
"00000000100001100100101110001010",
"00000000100001101001001000100010",
"00000000100001101101100100000101",
"00000000100001110010000000110010",
"00000000100001110110011110101011",
"00000000100001111010111101101111",
"00000000100001111111011110000000",
"00000000100010000011111111011101",
"00000000100010001000100010001000",
"00000000100010001101000110000000",
"00000000100010010001101011000111",
"00000000100010010110010001011100",
"00000000100010011010111001000000",
"00000000100010011111100001110100",
"00000000100010100100001011111000",
"00000000100010101000110111001101",
"00000000100010101101100011110010",
"00000000100010110010010001101010",
"00000000100010110111000000110100",
"00000000100010111011110001010000",
"00000000100011000000100011000000",
"00000000100011000101010110000100",
"00000000100011001010001010011100",
"00000000100011001111000000001000",
"00000000100011010011110111001011",
"00000000100011011000101111100011",
"00000000100011011101101001010010",
"00000000100011100010100100010111",
"00000000100011100111100000110101",
"00000000100011101100011110101011",
"00000000100011110001011101111001",
"00000000100011110110011110100001",
"00000000100011111011100000100011",
"00000000100100000000100100000000",
"00000000100100000101101000111000",
"00000000100100001010101111001100",
"00000000100100001111110110111100",
"00000000100100010101000000001001",
"00000000100100011010001010110011",
"00000000100100011111010110111100",
"00000000100100100100100100100100",
"00000000100100101001110011101011",
"00000000100100101111000100010011",
"00000000100100110100010110011011",
"00000000100100111001101010000101",
"00000000100100111110111111010001",
"00000000100101000100010110000000",
"00000000100101001001101110010010",
"00000000100101001111001000001001",
"00000000100101010100100011100100",
"00000000100101011010000000100101",
"00000000100101011111011111001100",
"00000000100101100100111111011010",
"00000000100101101010100001010000",
"00000000100101110000000100101110",
"00000000100101110101101001110101",
"00000000100101111011010000100101",
"00000000100110000000111001000001",
"00000000100110000110100011001000",
"00000000100110001100001110111010",
"00000000100110010001111100011010",
"00000000100110010111101011100111",
"00000000100110011101011100100010",
"00000000100110100011001111001101",
"00000000100110101001000011100111",
"00000000100110101110111001110010",
"00000000100110110100110001101111",
"00000000100110111010101011011110",
"00000000100111000000100111000000",
"00000000100111000110100100010110",
"00000000100111001100100011100001",
"00000000100111010010100100100001",
"00000000100111011000100111011000",
"00000000100111011110101100000110",
"00000000100111100100110010101101",
"00000000100111101010111011001100",
"00000000100111110001000101100101",
"00000000100111110111010001111010",
"00000000100111111101100000001001",
"00000000101000000011110000010110",
"00000000101000001010000010100000",
"00000000101000010000010110101001",
"00000000101000010110101100110001",
"00000000101000011101000100111001",
"00000000101000100011011111000011",
"00000000101000101001111011001111",
"00000000101000110000011001011110",
"00000000101000110110111001110001",
"00000000101000111101011100001010",
"00000000101001000100000000101001",
"00000000101001001010100111001111",
"00000000101001010001001111111101",
"00000000101001010111111010110101",
"00000000101001011110100111110110",
"00000000101001100101010111000100",
"00000000101001101100001000011101",
"00000000101001110010111100000101",
"00000000101001111001110001111011",
"00000000101010000000101010000000",
"00000000101010000111100100010111",
"00000000101010001110100000111111",
"00000000101010010101011111111010",
"00000000101010011100100001001010",
"00000000101010100011100100101111",
"00000000101010101010101010101010",
"00000000101010110001110010111101",
"00000000101010111000111101101001",
"00000000101011000000001010110000",
"00000000101011000111011010010001",
"00000000101011001110101100001111",
"00000000101011010110000000101011",
"00000000101011011101010111100110",
"00000000101011100100110001000001",
"00000000101011101100001100111110",
"00000000101011110011101011011101",
"00000000101011111011001100100001",
"00000000101100000010110000001011",
"00000000101100001010010110011011",
"00000000101100010001111111010011",
"00000000101100011001101010110101",
"00000000101100100001011001000010",
"00000000101100101001001001111100",
"00000000101100110000111101100011",
"00000000101100111000110011111001",
"00000000101101000000101101000000",
"00000000101101001000101000111001",
"00000000101101010000100111100110",
"00000000101101011000101001001000",
"00000000101101100000101101100000",
"00000000101101101000110100110001",
"00000000101101110000111110111011",
"00000000101101111001001100000000",
"00000000101110000001011100000010",
"00000000101110001001101111000011",
"00000000101110010010000101000011",
"00000000101110011010011110000110",
"00000000101110100010111010001011",
"00000000101110101011011001010110",
"00000000101110110011111011100111",
"00000000101110111100100001000000",
"00000000101111000101001001100100",
"00000000101111001101110101010011",
"00000000101111010110100100010000",
"00000000101111011111010110011100",
"00000000101111101000001011111010",
"00000000101111110001000100101010",
"00000000101111111010000000101111",
"00000000110000000011000000001100",
"00000000110000001100000011000000",
"00000000110000010101001001010000",
"00000000110000011110010010111011",
"00000000110000100111100000000110",
"00000000110000110000110000110000",
"00000000110000111010000100111101",
"00000000110001000011011100101111",
"00000000110001001100111000000111",
"00000000110001010110010111001000",
"00000000110001011111111001110100",
"00000000110001101001100000001100",
"00000000110001110011001010010011",
"00000000110001111100111000001100",
"00000000110010000110101001111000",
"00000000110010010000011111011010",
"00000000110010011010011000110011",
"00000000110010100100010110000111",
"00000000110010101110010111011000",
"00000000110010111000011100100111",
"00000000110011000010100101111000",
"00000000110011001100110011001100",
"00000000110011010111000100100111",
"00000000110011100001011010001010",
"00000000110011101011110011111000",
"00000000110011110110010001110100",
"00000000110100000000110100000000",
"00000000110100001011011010011111",
"00000000110100010110000101010100",
"00000000110100100000110100100000",
"00000000110100101011101000001000",
"00000000110100110110100000001101",
"00000000110101000001011100110010",
"00000000110101001100011101111011",
"00000000110101010111100011101001",
"00000000110101100010101110000000",
"00000000110101101101111101000011",
"00000000110101111001010000110101",
"00000000110110000100101001011001",
"00000000110110010000000110110010",
"00000000110110011011101001000010",
"00000000110110100111010000001101",
"00000000110110110010111100010111",
"00000000110110111110101101100001",
"00000000110111001010100011110001",
"00000000110111010110011111001000",
"00000000110111100010011111101011",
"00000000110111101110100101011100",
"00000000110111111010110000011111",
"00000000111000000111000000111000",
"00000000111000010011010110101001",
"00000000111000011111110001111000",
"00000000111000101100010010100110",
"00000000111000111000111000111000",
"00000000111001000101100100110010",
"00000000111001010010010110011000",
"00000000111001011111001101101100",
"00000000111001101100001010110100",
"00000000111001111001001101110010",
"00000000111010000110010110101100",
"00000000111010010011100101100101",
"00000000111010100000111010100000",
"00000000111010101110010101100100",
"00000000111010111011110110110010",
"00000000111011001001011110010001",
"00000000111011010111001100000011",
"00000000111011100101000000001110",
"00000000111011110010111010110111",
"00000000111100000000111100000000",
"00000000111100001111000011110000",
"00000000111100011101010010001011",
"00000000111100101011100111010110",
"00000000111100111010000011010101",
"00000000111101001000100110001101",
"00000000111101010111010000000011",
"00000000111101100110000000111101",
"00000000111101110100111000111111",
"00000000111110000011111000001111",
"00000000111110010010111110110010",
"00000000111110100010001100101100",
"00000000111110110001100010000101",
"00000000111111000000111111000000",
"00000000111111010000100011100101",
"00000000111111100000001111111000",
"00000000111111110000000011111111",
"00000001000000000000000000000000",
"00000001000000010000000100000001",
"00000001000000100000010000001000",
"00000001000000110000100100011011",
"00000001000001000001000001000001",
"00000001000001010001100101111111",
"00000001000001100010010011011101",
"00000001000001110011001001100000",
"00000001000010000100001000010000",
"00000001000010010101001111110011",
"00000001000010100110100000010000",
"00000001000010110111111001101110",
"00000001000011001001011100010100",
"00000001000011011011001000001010",
"00000001000011101100111101010110",
"00000001000011111110111100000001",
"00000001000100010001000100010001",
"00000001000100100011010110001110",
"00000001000100110101110010000001",
"00000001000101001000010111110000",
"00000001000101011011000111100101",
"00000001000101101110000001101000",
"00000001000110000001000110000001",
"00000001000110010100010100111000",
"00000001000110100111101110010110",
"00000001000110111011010010100100",
"00000001000111001111000001101010",
"00000001000111100010111011110011",
"00000001000111110111000001000111",
"00000001001000001011010001110000",
"00000001001000011111101101111000",
"00000001001000110100010101100111",
"00000001001001001001001001001001",
"00000001001001011110001000100111",
"00000001001001110011010100001011",
"00000001001010001000101100000001",
"00000001001010011110010000010010",
"00000001001010110100000001001010",
"00000001001011001001111110110100",
"00000001001011100000001001011100",
"00000001001011110110100001001011",
"00000001001100001101000110010000",
"00000001001100100011111000110100",
"00000001001100111010111001000101",
"00000001001101010010000111001111",
"00000001001101101001100011011111",
"00000001001110000001001110000001",
"00000001001110011001000111000010",
"00000001001110110001001110110001",
"00000001001111001001100101011010",
"00000001001111100010001011001011",
"00000001001111111011000000010011",
"00000001010000010100000101000001",
"00000001010000101101011001100010",
"00000001010001000110111110000110",
"00000001010001100000110010111100",
"00000001010001111010111000010100",
"00000001010010010101001110011110",
"00000001010010101111110101101010",
"00000001010011001010101110001000",
"00000001010011100101111000001010",
"00000001010100000001010100000001",
"00000001010100011101000001111110",
"00000001010100111001000010010100",
"00000001010101010101010101010101",
"00000001010101110001111011010011",
"00000001010110001110110100100011",
"00000001010110101100000001010110",
"00000001010111001001100010000010",
"00000001010111100111010110111011",
"00000001011000000101100000010110",
"00000001011000100011111110100111",
"00000001011001000010110010000101",
"00000001011001100001111011000110",
"00000001011010000001011010000001",
"00000001011010100001001111001101",
"00000001011011000001011011000001",
"00000001011011100001111101110110",
"00000001011100000010111000000101",
"00000001011100100100001010000111",
"00000001011101000101110100010111",
"00000001011101100111110111001110",
"00000001011110001010010011001000",
"00000001011110101101001000100000",
"00000001011111010000010111110100",
"00000001011111110100000001011111",
"00000001100000011000000110000001",
"00000001100000111100100101110111",
"00000001100001100001100001100001",
"00000001100010000110111001011111",
"00000001100010101100101110010000",
"00000001100011010011000000011000",
"00000001100011111001110000011000",
"00000001100100100000111110110100",
"00000001100101001000101100001111",
"00000001100101110000111001001111",
"00000001100110011001100110011001",
"00000001100111000010110100010100",
"00000001100111101100100011101001",
"00000001101000010110110100111111",
"00000001101001000001101001000001",
"00000001101001101101000000011010",
"00000001101010011000111011110110",
"00000001101011000101011100000001",
"00000001101011110010100001101011",
"00000001101100100000001101100100",
"00000001101101001110100000011011",
"00000001101101111101011011000011",
"00000001101110101100111110010001",
"00000001101111011101001010111000",
"00000001110000001110000001110000",
"00000001110000111111100011110000",
"00000001110001110001110001110001",
"00000001110010100100101100110000",
"00000001110011011000010101101000",
"00000001110100001100101101011000",
"00000001110101000001110101000001",
"00000001110101110111101101100101",
"00000001110110101110011000000111",
"00000001110111100101110101101110",
"00000001111000011110000111100001",
"00000001111001010111001110101100",
"00000001111010010001001100011010",
"00000001111011001100000001111011",
"00000001111100000111110000011111",
"00000001111101000100011001011001",
"00000001111110000001111110000001",
"00000001111111000000011111110000",
"00000010000000000000000000000000",
"00000010000001000000100000010000",
"00000010000010000010000010000010",
"00000010000011000100100110111010",
"00000010000100001000010000100001",
"00000010000101001101000000100001",
"00000010000110010010111000101001",
"00000010000111011001111010101101",
"00000010001000100010001000100010",
"00000010001001101011100100000010",
"00000010001010110110001111001011",
"00000010001100000010001100000010",
"00000010001101001111011100101100",
"00000010001110011110000011010101",
"00000010001111101110000010001111",
"00000010010000111111011011110000",
"00000010010010010010010010010010",
"00000010010011100110101000010111",
"00000010010100111100100000100101",
"00000010010110010011111101101001",
"00000010010111101101000010010111",
"00000010011001000111110001101001",
"00000010011010100100001110011111",
"00000010011100000010011100000010",
"00000010011101100010011101100010",
"00000010011111000100010110010111",
"00000010100000101000001010000010",
"00000010100010001101111100001100",
"00000010100011110101110000101000",
"00000010100101011111101011010100",
"00000010100111001011110000010100",
"00000010101000111010000011111101",
"00000010101010101010101010101010",
"00000010101100011101101001000110",
"00000010101110010011000100000101",
"00000010110000001011000000101100",
"00000010110010000101100100001011",
"00000010110100000010110100000010",
"00000010110110000010110110000010",
"00000010111000000101110000001011",
"00000010111010001011101000101110",
"00000010111100010100100110010000",
"00000010111110100000101111101000",
"00000011000000110000001100000011",
"00000011000011000011000011000011",
"00000011000101011001011100100001",
"00000011000111110011100000110001",
"00000011001010010001011000011111",
"00000011001100110011001100110011",
"00000011001111011001000111010010",
"00000011010010000011010010000011",
"00000011010100110001110111101100",
"00000011010111100101000011010111",
"00000011011010011101000000110110",
"00000011011101011001111100100010",
"00000011100000011100000011100000",
"00000011100011100011100011100011",
"00000011100110110000101011010001",
"00000011101010000011101010000011",
"00000011101101011100110000001110",
"00000011110000111100001111000011",
"00000011110100100010011000110101",
"00000011111000001111100000111110",
"00000011111100000011111100000011",
"00000100000000000000000000000000",
"00000100000100000100000100000100",
"00000100001000010000100001000010",
"00000100001100100101110001010011",
"00000100010001000100010001000100",
"00000100010101101100011110010111",
"00000100011010011110111001011000",
"00000100011111011100000100011111",
"00000100100100100100100100100100",
"00000100101001111001000001001010",
"00000100101111011010000100101111",
"00000100110101001000011100111110",
"00000100111011000100111011000100",
"00000101000001010000010100000101",
"00000101000111101011100001010001",
"00000101001110010111100000101001",
"00000101010101010101010101010101",
"00000101011100100110001000001010",
"00000101100100001011001000010110",
"00000101101100000101101100000101",
"00000101110100010111010001011101",
"00000101111101000001011111010000",
"00000110000110000110000110000110",
"00000110001111100111000001100011",
"00000110011001100110011001100110",
"00000110100100000110100100000110",
"00000110101111001010000110101111",
"00000110111010110011111001000101",
"00000111000111000111000111000111",
"00000111010100000111010100000111",
"00000111100001111000011110000111",
"00000111110000011111000001111100",
"00001000000000000000000000000000",
"00001000010000100001000010000100",
"00001000100010001000100010001000",
"00001000110100111101110010110000",
"00001001001001001001001001001001",
"00001001011110110100001001011110",
"00001001110110001001110110001001",
"00001010001111010111000010100011",
"00001010101010101010101010101010",
"00001011001000010110010000101100",
"00001011101000101110100010111010",
"00001100001100001100001100001100",
"00001100110011001100110011001100",
"00001101011110010100001101011110",
"00001110001110001110001110001110",
"00001111000011110000111100001111",
"00010000000000000000000000000000",
"00010001000100010001000100010001",
"00010010010010010010010010010010",
"00010011101100010011101100010011",
"00010101010101010101010101010101",
"00010111010001011101000101110100",
"00011001100110011001100110011001",
"00011100011100011100011100011100",
"00100000000000000000000000000000",
"00100100100100100100100100100100",
"00101010101010101010101010101010",
"00110011001100110011001100110011",
"01000000000000000000000000000000",
"01010101010101010101010101010101",
"10000000000000000000000000000000"
 );
begin

INIT : process(DENOMINATOR,RESET)
begin
	if RESET = '1' then
		DENOMINATOR2 <= "0000000010";
	else
		DENOMINATOR2 <= DENOMINATOR;
	end if;
end process INIT;

SETNUMERATOR : process (CLOCK)
begin
	if CLOCK'event and CLOCK = '1' then
		if RESET = '1' then
			NUMERATOR2 <= "0000000001";
		else
			NUMERATOR2 <= NUMERATOR;
		end if;
	end if;
end process SETNUMERATOR;
			

INDEX <= DENOMINATOR2 - "0000000010";

LOOKUP: process(CLOCK)
begin
	if CLOCK'event and CLOCK = '1' then
		 RECIPROCAL <= LUT(conv_integer(INDEX));
	end if;
end process LOOKUP;

DIVIDE1: process(CLOCK)
begin
	if CLOCK'event and CLOCK='1' then
		PRODUCT1<=NUMERATOR2*RECIPROCAL(31 downto 16);
	end if;
end process DIVIDE1;

DIVIDE2: process(CLOCK)
begin
	if CLOCK'event and CLOCK='1' then
		PRODUCT2<=NUMERATOR2*RECIPROCAL(15 downto 0);
	end if;
end process DIVIDE2;

TOTAL<=((PRODUCT1 & "0000000000000000") + ("0000000000000000" & PRODUCT2));
QUOTIENT <=	 TOTAL(31 downto 22);


end RTL;
